library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
	
package port_dizi_paket is
	
  type port_dizi is array (3 downto 0) of std_logic_vector(0 to 7);

end port_dizi_paket;